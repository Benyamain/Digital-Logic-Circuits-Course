`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02/22/2024 05:18:46 PM
// Design Name: 
// Module Name: 1bit_full_adder_3
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module 1bit_full_adder_3(
    input a,
    input b,
    input cin,
    output s,
    output cout
    );
endmodule
